	component oscillator is
		port (
			oscena : in  std_logic := 'X'; -- oscena
			clkout : out std_logic         -- clkout
		);
	end component oscillator;

	u0 : component oscillator
		port map (
			oscena => CONNECTED_TO_oscena, -- oscena.oscena
			clkout => CONNECTED_TO_clkout  -- clkout.clkout
		);

