
module clock_100ms (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
