// clock_100ms.v

// Generated using ACDS version 14.0 200 at 2014.11.30.16:36:37

`timescale 1 ps / 1 ps
module clock_100ms (
		input  wire  inclk,  //  altclkctrl_input.inclk
		output wire  outclk  // altclkctrl_output.outclk
	);

	clock_100ms_altclkctrl_0 altclkctrl_0 (
		.inclk  (inclk),  //  altclkctrl_input.inclk
		.outclk (outclk)  // altclkctrl_output.outclk
	);

endmodule
